module timeset()
